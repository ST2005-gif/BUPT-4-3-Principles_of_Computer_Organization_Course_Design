module ver2 (
        //����˿�
        input wire [2:0] SWC_SWB_SWA,      // ģʽѡ���ź�
        input wire [3:0] IR7_IR4
,          // ָ��Ĵ�����4λ
        input wire CLR,                    // ��λ�ź� (����Ч)
        input wire T3,                     // ʱ���ź� T3 (��ΪST0��ʱ��)
        input wire W1, W2, W3,             // ΢ָ��ʱ���ź�
        input wire C, Z,                   // ״̬��־����λC����Z
        //����˿�
        output reg SELCTL,                 // ѡ������ź�
        output reg ABUS,                   // ����ALU�����Ƿ������������
        output reg SBUS,                   // �����ֶ����������Ƿ������������
        output reg MBUS,                   // ����˫�˿ڴ洢���������͵���������
        output reg M,CIN,                  // M�ǿ���ALU���߼����㻹���������� CIN��������S���M��Ӧ�Ĳ������н�λ���������޽�λ����
        output reg DRW,                    // ���ƼĴ���д���ź�
        output reg LDZ,                    // ��Ϊ1����������Ϊ0ʱ��ZΪ1������Ϊ0����ZΪ0
        output reg LDC,                    // ��Ϊ1����������������λʱ��CΪ1�����޽�λ����CΪ0
        output reg MEMW,                   // ���ƴ洢��˫�˿�RAMд���źţ�Ϊ1ʱ�������е�ֵд�봢����
        output reg ARINC,                  // ���Ƶ�ַ�Ĵ���AR��ֵ��1�ź�
        output reg PCINC,                  // ���Ƶ�ַ�Ĵ���PC��ֵ��1�ź�
        output reg PCADD,                  // ����PC��ָ���ַ�ź�
        output reg LPC,                    // ���ƽ���������������д��PC�Ĵ���
        output reg LAR,                    // ���ƽ���������������д��AR�Ĵ���
        output reg LIR,                    // ���ƽ���������������д��IR�Ĵ���
        output reg STOP,                   // ֹͣ�ź�
        output reg SHORT,                  // ����ʱ�ź�
        output reg LONG,                   // ����ʱ�ź�
        output reg [3:0] S, SEL            // S����ALU������ͬ�ĺ��� SEL���� 2 - 4 ������
    );
    //״̬��ʶ
    // �ڲ��ź�����
    reg ST0;
    wire WRITE_REG, READ_REG, INS_FETCH, WRITE_MEM, READ_MEM;
    wire ADD, SUB, AND, INC, LD, ST, JC, JZ, JMP, STP;
    wire NOP, OUT, NOT, CMP, MOV, DEC;
    reg [3:1] W; // ���ڴ洢W�źŵ�״̬
    wire short_command;
    wire long_command;

    // �ڽ���׶�ȷ��ָ���
    assign short_command = (NOP || ADD || SUB || AND || INC || (JC && !C) ||
                         (JZ && !Z) || OUT || NOT || CMP || MOV || DEC ||
                         READ_MEM || WRITE_MEM);

    assign long_command = 1'b0;

    // T3�½��ؼ������߼�
    always @(negedge T3 or negedge CLR) begin
        if (!CLR) begin
            W[1] <= 1'b1;
            W[2] <= 1'b0;
            W[3] <= 1'b0;
        end
        else begin
            if(W[1]) begin
                if(short_command) begin
                    W[1] <= 1'b1;
                    W[2] <= 1'b0;
                    W[3] <= 1'b0;
                end
                else begin
                    W[1] <= 1'b0;
                    W[2] <= 1'b1;
                    W[3] <= 1'b0;
                end
            end
            else if(W[2]) begin
                if(long_command) begin
                    W[1] <= 1'b0;
                    W[2] <= 1'b0;
                    W[3] <= 1'b1;
                end
                else begin
                    W[1] <= 1'b1;
                    W[2] <= 1'b0;
                    W[3] <= 1'b0;
                end
            end
            else if(W[3]) begin
                W[1] <= 1'b1;
                W[2] <= 1'b0;
                W[3] <= 1'b0; // ����Ϊ��ʼ״̬
            end
        end
    end

    // ST0״̬�� - ָ��ִ��״̬
    always @(negedge T3 or negedge CLR) begin
        if (!CLR) begin
            ST0 <= 1'b0;
        end
        else begin
            if (!ST0 && ((WRITE_REG && W[2]) || (READ_MEM && W[1]) ||
                         (WRITE_MEM && W[1]) || (INS_FETCH && W[2]))) begin
                ST0 <= 1'b1;
            end
            else if (ST0 && (WRITE_REG && W[2])) begin
                ST0 <= 1'b0;
            end
        end
    end

    // ����ģʽ����
    assign WRITE_REG = (SWC_SWB_SWA == 3'b100);
    assign READ_REG = (SWC_SWB_SWA == 3'b011);
    assign INS_FETCH = (SWC_SWB_SWA == 3'b000);
    assign READ_MEM = (SWC_SWB_SWA == 3'b010);
    assign WRITE_MEM = (SWC_SWB_SWA == 3'b001);

    // ָ������
    assign ADD = (IR7_IR4 == 4'b0001) && INS_FETCH && ST0;
    assign SUB = (IR7_IR4 == 4'b0010) && INS_FETCH && ST0;
    assign AND = (IR7_IR4 == 4'b0011) && INS_FETCH && ST0;
    assign INC = (IR7_IR4 == 4'b0100) && INS_FETCH && ST0;
    assign LD = (IR7_IR4 == 4'b0101) && INS_FETCH && ST0;
    assign ST = (IR7_IR4 == 4'b0110) && INS_FETCH && ST0;
    assign JC = (IR7_IR4 == 4'b0111) && INS_FETCH && ST0;
    assign JZ = (IR7_IR4 == 4'b1000) && INS_FETCH && ST0;
    assign JMP = (IR7_IR4 == 4'b1001) && INS_FETCH && ST0;
    assign STP = (IR7_IR4 == 4'b1110) && INS_FETCH && ST0;
    assign NOP = (IR7_IR4 == 4'b0000) && INS_FETCH && ST0;
    assign OUT = (IR7_IR4 == 4'b1010) && INS_FETCH && ST0;
    assign NOT = (IR7_IR4 == 4'b1101) && INS_FETCH && ST0;
    assign CMP = (IR7_IR4 == 4'b1100) && INS_FETCH && ST0;
    assign MOV = (IR7_IR4 == 4'b1011) && INS_FETCH && ST0;
    assign DEC = (IR7_IR4 == 4'b1111) && INS_FETCH && ST0;

    // ȫʱ���߼����� - ���п����ź���T3�½��ظ���
    always @(negedge T3 or negedge CLR) begin
        if (!CLR) begin
            // ��λ���п����ź�
            SELCTL <= 1'b0;
            DRW <= 1'b0;
            LPC <= 1'b0;
            PCINC <= 1'b0;
            PCADD <= 1'b0;
            LAR <= 1'b0;
            ARINC <= 1'b0;
            LIR <= 1'b0;
            LDZ <= 1'b0;
            LDC <= 1'b0;
            CIN <= 1'b0;
            M <= 1'b0;
            MEMW <= 1'b0;
            ABUS <= 1'b0;
            SBUS <= 1'b0;
            MBUS <= 1'b0;
            STOP <= 1'b0;
            SHORT <= 1'b0;
            LONG <= 1'b0;
            S <= 4'b0000;
            SEL <= 4'b0000;
        end
        else begin
            // �����źźϳ� - ���п����ź�ͬ������
            SBUS <= (WRITE_REG && (W[1] || W[2])) || (READ_MEM && (W[1] && !ST0)) ||
                 (WRITE_MEM && W[1]) || (INS_FETCH && (W[1] && !ST0));

            SEL[3] <= (WRITE_REG && (W[1] || W[2]) && ST0) || (READ_REG && W[2]);
            SEL[2] <= WRITE_REG && W[2];
            SEL[1] <= (WRITE_REG && ((W[1] && !ST0) || (W[2] && ST0))) || (READ_REG && W[2]);
            SEL[0] <= (WRITE_REG && W[1]) || (READ_REG && (W[1] || W[2]));

            SELCTL <= ((WRITE_REG || READ_REG) && (W[1] || W[2])) || ((READ_MEM || WRITE_MEM) && W[1]);

            DRW <= (WRITE_REG && (W[1] || W[2])) ||
                ((ADD || SUB || AND || INC || NOT || MOV || DEC) && W[1]) ||
                (LD && W[2]);

            STOP <= ((WRITE_REG || READ_REG) && (W[1] || W[2])) ||
                 ((READ_MEM || WRITE_MEM) && W[1]) ||
                 (STP && W[1]) ||
                 (INS_FETCH && !ST0 && W[1]);

            LAR <= ((READ_MEM || WRITE_MEM) && W[1] && !ST0) || ((ST || LD) && W[1]);

            SHORT <= ((READ_MEM || WRITE_MEM) && W[1]) ||
                  ((NOP || ADD || SUB || AND || INC || (JC && !C) ||
                    (JZ && !Z) || OUT || NOT || CMP || MOV) && W[1]);

            MBUS <= (READ_MEM && W[1] && ST0) || (LD && W[2]);

            ARINC <= (WRITE_MEM || READ_MEM) && W[1] && ST0;

            MEMW <= (WRITE_MEM && W[1] && ST0) || (ST && W[2]);

            CIN <= (ADD || DEC)&& W[1];

            ABUS <= ((ADD || SUB || AND || INC || LD || ST || JMP || OUT || MOV || CMP || NOT || DEC) && W[1]) ||
                 (ST && W[2]);

            LDZ <= (ADD || SUB || AND || INC || CMP || DEC) && W[1];
            LDC <= (ADD || SUB || INC || CMP || NOT || DEC) && W[1];

            M <= ((AND || LD || ST || JMP || OUT || MOV || NOT) && W[1]) ||
              (ST && W[2]);

            S[3] <= ((ADD || AND || LD || ST || JMP || OUT || MOV || DEC) && W[1]) ||
             (ST && W[2]);
            S[2] <= ((SUB || ST || JMP || CMP || DEC) && W[1]);
            S[1] <= ((SUB || AND || LD || ST || JMP || OUT || MOV || CMP || DEC) && W[1]) ||
             (ST && W[2]);
            S[0] <= (ADD || AND || ST || JMP || DEC) && W[1];

            LPC <= (JMP && W[1]) || (INS_FETCH && !ST0 && W[1]);

            LONG <= 1'b0; // û�����ó����ڿ���

            PCADD <= ((C && JC) || (Z && JZ)) && W[1];

            // �ȸ���LIR�ź�
            LIR <= (INS_FETCH && W[2] && !ST0) ||
                ((NOP || ADD || SUB || AND || INC || (JC && !C) ||
                  (JZ && !Z) || OUT || MOV || CMP || NOT) && W[1]) ||
                ((LD || ST || (JC && C) || (JZ && Z) || JMP) && W[2]);

            // �����PCINC�ź�
            PCINC <= (INS_FETCH && W[2] && !ST0) ||
                  ((NOP || ADD || SUB || AND || INC || (JC && !C) ||
                    (JZ && !Z) || OUT || MOV || CMP || NOT) && W[1]) ||
                  ((LD || ST || (JC && C) || (JZ && Z) || JMP) && W[2]);
        end
    end

endmodule

